`ifndef _CPU_PARAM_SV 
`define _CPU_PARAM_SV
package cpu_param;










endpackage
`endif 


