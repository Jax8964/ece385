`ifndef _CONST_SV
`define _CONST_SV

`define CLOCK_PERIOD    24
`define FLAG_N SR[7]
`define FLAG_V SR[6]
`define FLAG_D SR[3]
`define FLAG_I SR[2]
`define FLAG_Z SR[1]
`define FLAG_C SR[0]

`define PPU_PERIOD    8




`endif
